
library IEEE;
use IEEE.STD_LOGIC_1164.all;

package Cards_Constants is
	
	constant Card_X	: integer := 66;
	constant Card_Y	: integer := 100;

	constant Numbers_Block_X	: integer := 16;
	constant Numbers_Block_Y	: integer := 16;
	
	constant Numbers_Block_X_0	: integer := 15;
	constant Numbers_Block_Y_0	: integer := 15;
	
	constant Numbers_Block_Size_0	: integer := 255;
	constant Numbers_Block_Size	: integer := 256;

	constant Numbers_Total_Size	: integer := 6656;
	constant Numbers_Total_Size_0	: integer := 6655;


	constant Seeds_Block_X	: integer := 32;
	constant Seeds_Block_X_0	: integer := 31;
	
	constant Seeds_Block_Y	: integer := 32;	
	constant Seeds_Block_Y_0	: integer := 31;

	constant Seeds_Block_Size	: integer := 1024;
	constant Seeds_Block_Size_0	: integer := 1023;

	constant Seeds_Total_Size	: integer := 4096;
	constant Seeds_Total_Size_0	: integer := 4095;


	constant Card_1_X : integer := 14;
	constant Card_1_Y : integer := 15;
	constant Card_2_X : integer := 94;
	constant Card_2_Y : integer := 15;
	constant Card_3_X : integer := 174;
	constant Card_3_Y : integer := 15;
	constant Card_4_X : integer := 14;
	constant Card_4_Y : integer := 130;
	constant Card_5_X : integer := 94;
	constant Card_5_Y : integer := 130;

	constant Card_D_1_X : integer := 14;
	constant Card_D_1_Y : integer := 15;
	constant Card_D_2_X : integer := 94;
	constant Card_D_2_Y : integer := 15;
	constant Card_D_3_X : integer := 174;
	constant Card_D_3_Y : integer := 15;
	constant Card_D_4_X : integer := 254;
	constant Card_D_4_Y : integer := 15;
	constant Card_D_5_X : integer := 334;
	constant Card_D_5_Y : integer := 15;

end Cards_Constants;

package body Cards_Constants is
 
end Cards_Constants;




	--constant Asso 			: integer := 0;
	--constant Asso_Red 		: integer := 256;
	--constant Due 			: integer := 512;
	--constant Due_Red 		: integer := 768;
	--constant Tre 			: integer := 1024;
	--constant Tre_Red 		: integer := 1280;
	--constant Quattro		: integer := 1536;
	--constant Quattro_Red 	: integer := 1792;
	--constant Cinque 		: integer := 2048;
	--constant Cinque_Red 	: integer := 2304;
	--constant Sei	 		: integer := 2560;
	--constant Sei_Red		: integer := 2816;
	--constant Sette	 		: integer := 3072;
	--constant Sette_Red	 	: integer := 3328;
	--constant Otto	 		: integer := 3584;
	--constant Otto_Red	 	: integer := 3840;
	--constant Nove 			: integer := 4096;
	--constant Nove_Red 		: integer := 4352;
	--constant Dieci			: integer := 4608;
	--constant Dieci_Red 		: integer := 4864;
	--constant Jack			: integer := 5120;
	--constant Jack_Red	 	: integer := 5376;
	--constant Queen	 		: integer := 5632;
	--constant Queen_Red 		: integer := 5888;
	--constant King	 		: integer := 6144;
	--constant King_Red 		: integer := 6400;
